/*
 this module implements bitwise OR operation for 32 bit vectors
 assign out = inA | inB;
 */
module bitwise_or (input [31:0] inA,
                   input [31:0] inB,
                   output [31:0] out);
assign out = 32'h00000000;
endmodule
